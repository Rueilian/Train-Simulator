module Time_display (
    input i_en,
    input i_minus,
    input [12:0] i_H_Cont,
    input [12:0] i_V_Cont,
    input [12:0] i_x,
    input [12:0] i_y,
    input [3:0] i_time,
    output reg o_valid
);

parameter WIDTH = 18;
parameter HEIGHT = 25;

wire [WIDTH*HEIGHT-1:0] number[0:9];
wire [WIDTH*HEIGHT-1:0] minus;
reg [WIDTH*HEIGHT-1:0] index;

assign number[0] = 450'b000000000000000000000000000000000000000000000000000000000000001111000000000000111111100000000001110001110000000011100000110000000011000000011000000010000000011000000110000000001000000110000000001100000110000000001100000110000000001000000100000000011000001100000000011000001100000000011000001100000000011000001100000000011000001100000000110000000110000001110000000111000011100000000011111111000000000000111100000000000000000000000000000000000000000000;
assign number[1] = 450'b000000000000000000000000000000000000000000000000000000000000000110000000000000001110000000000000011110000000000000000110000000000000000110000000000000001100000000000000001100000000000000001100000000000000001100000000000000001100000000000000001100000000000000001100000000000000001100000000000000001100000000000000011000000000000000011000000000000000011000000000000000011000000000000000010000000000000000000000000000000000000000000000000000000000000000;
assign number[2] = 450'b000000000000000000000000000000000000000000000000000000000000011111100000000001111111110000000011100000111000000011000000011000000110000000001100000110000000001100000000000000001100000000000000011000000000000000111000000000000001110000000000011111100000000001111110000000000011100000000000000110000000000000000110000000000000001100000000000000001100000000000000001111111111110000001111111111111000000000000000000000000000000000000000000000000000000000;
assign number[3] = 450'b000000000000000000000000000000000000000000000000000000000000011111000000000000111111100000000000110001110000000000000000110000000000000000110000000000000000110000000000000011100000000000000111000000000000000111100000000000000001110000000000000000011000000000000000011000000000000000011000000000000000011000000000000000011000000110000000110000000111000011110000000011111111100000000001111110000000000000000000000000000000000000000000000000000000000000;
assign number[4] = 450'b000000000000000000000000000000000000000000000000000000000000000001100000000000000011110000000000000011110000000000000110110000000000000110100000000000001100100000000000001101100000000000011001100000000000011001100000000000110011000000000001100011000000000011111111111000000111111111111000000000000011000000000000000011000000000000000011000000000000000011000000000000000010000000000000000010000000000000000000000000000000000000000000000000000000000000;
assign number[5] = 450'b000000000000000000000000000000000000000000000000000000000001111111111000000001111111110000000001100000000000000001100000000000000001100000000000000011000000000000000011000000000000000011111111000000000011111111100000000000000001110000000000000000110000000000000000011000000000000000011000001100000000011000001100000000011000000110000000110000000111000001110000000011111111100000000001111110000000000000000000000000000000000000000000000000000000000000;
assign number[6] = 450'b000000000000000000000000000000000000000000000000000000000000001110000000000000111111100000000001110001110000000011000000000000000011000000000000000110000000000000000110000000000000000110001110000000000110111111100000000111110001110000001111000000110000001110000000111000001100000000011000001100000000011000001100000000011000001100000000110000000110000001110000000111000011100000000011111111000000000000111110000000000000000000000000000000000000000000;
assign number[7] = 450'b000000000000000000000000000000000000000000000000000000001111111111111100000111111111111100000000000000011000000000000000110000000000000001100000000000000001100000000000000011000000000000000110000000000000000110000000000000001100000000000000011000000000000000011000000000000000110000000000000001100000000000000001100000000000000011000000000000000110000000000000000110000000000000001100000000000000001000000000000000000000000000000000000000000000000000;
assign number[8] = 450'b000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000111001100000000001110000110000000001100000110000000001100000110000000001100001100000000000110011100000000000111111000000000001110011100000000011000000110000000110000000011000000110000000011000001100000000011000001100000000011000001110000000010000000110000000110000000111000011100000000011111111000000000001111110000000000000000000000000000000000000000000;
assign number[9] = 450'b000000000000000000000000000000000000000000000000000000000000001111000000000000111111110000000001110001110000000011100000011000000011000000011000000110000000001100000110000000001100000110000000001100000110000000011000000011000000111000000011100011111000000001111111011000000000011100011000000000000000011000000000000000011000000000000000110000000000000001110000000011000011100000000011111111000000000000111100000000000000000000000000000000000000000000;
assign minus = 450'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000011111111111000000111111110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

always @(*) begin

    index = (WIDTH*HEIGHT - ( (i_V_Cont-i_y)*WIDTH+(i_H_Cont-i_x)+1 ));

    // valid
    if (i_en && i_H_Cont-i_x >= 0 && i_H_Cont-i_x < WIDTH && i_V_Cont-i_y >= 0 && i_V_Cont-i_y < HEIGHT) begin
        if (i_minus == 0) begin
            case (i_time)
                4'd0: begin o_valid = number[0][index]; end
                4'd1: begin o_valid = number[1][index]; end
                4'd2: begin o_valid = number[2][index]; end
                4'd3: begin o_valid = number[3][index]; end
                4'd4: begin o_valid = number[4][index]; end
                4'd5: begin o_valid = number[5][index]; end
                4'd6: begin o_valid = number[6][index]; end
                4'd7: begin o_valid = number[7][index]; end
                4'd8: begin o_valid = number[8][index]; end
                4'd9: begin o_valid = number[9][index]; end
                default: begin o_valid = 0; end
            endcase
        end else begin
            o_valid = minus[index];
        end
    end else begin
        o_valid = 0;
    end
end

endmodule