module Minus_display (
    input i_en,
    input [12:0] i_H_Cont,
    input [12:0] i_V_Cont,
    input [12:0] i_x,
    input [12:0] i_y,
    output reg o_valid
);

parameter WIDTH = 18;
parameter HEIGHT = 25;

wire [WIDTH*HEIGHT-1:0] minus;
reg [WIDTH*HEIGHT-1:0] index;

assign minus = 450'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000011111111111000000111111110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

always @(*) begin

    index = (WIDTH*HEIGHT - ( (i_V_Cont-i_y)*WIDTH+(i_H_Cont-i_x)+1 ));

    // valid
    if (i_en && i_H_Cont-i_x >= 0 && i_H_Cont-i_x < WIDTH && i_V_Cont-i_y >= 0 && i_V_Cont-i_y < HEIGHT) begin
        o_valid = minus[index];
    end else begin
        o_valid = 0;
    end
end

endmodule