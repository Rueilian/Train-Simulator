module Speed_display (
    input i_en,
    input [12:0] i_H_Cont,
    input [12:0] i_V_Cont,
    input [12:0] i_x,
    input [12:0] i_y,
    input [3:0] i_speed,
    output reg o_valid
);

parameter WIDTH = 18;
parameter HEIGHT = 30;

wire [WIDTH*HEIGHT-1:0] number[0:9];
reg [WIDTH*HEIGHT-1:0] index;

assign number[0] = 540'b000000000000000000_000000111111000000_000001111111100000_000100111111001000_001110000000011100_001111000000111100_001111000000111100_001111000000111100_001111000000111100_001111000000111100_001111000000111100_001111000000111100_001110000000011100_000100000000001000_000000000000000000_000100000000001000_001110000000011100_001111000000111100_001111000000111100_001111000000111100_001111000000111100_001111000000111100_001111000000111100_001111000000111100_001110000000011100_000100111111001000_000001111111100000_000000111111000000_000000000000000000_000000000000000000;
assign number[1] = 540'b000000000000000000_000000000000000000_000000000000000000_000000000000001000_000000000000011100_000000000000111100_000000000000111100_000000000000111100_000000000000111100_000000000000111100_000000000000111100_000000000000111100_000000000000011100_000000000000001000_000000000000000000_000000000000001000_000000000000011100_000000000000111100_000000000000111100_000000000000111100_000000000000111100_000000000000111100_000000000000111100_000000000000111100_000000000000011100_000000000000001000_000000000000000000_000000000000000000_000000000000000000_000000000000000000;
assign number[2] = 540'b000000000000000000_000000111111000000_000001111111100000_000000111111001000_000000000000011100_000000000000111100_000000000000111100_000000000000111100_000000000000111100_000000000000111100_000000000000111100_000000000000111100_000000000000011100_000000111111001000_000001111111100000_000100111111000000_001110000000000000_001111000000000000_001111000000000000_001111000000000000_001111000000000000_001111000000000000_001111000000000000_001111000000000000_001110000000000000_000100111111000000_000001111111100000_000000111111000000_000000000000000000_000000000000000000;
assign number[3] = 540'b000000000000000000_000000111111000000_000001111111100000_000000111111001000_000000000000011100_000000000000111100_000000000000111100_000000000000111100_000000000000111100_000000000000111100_000000000000111100_000000000000111100_000000000000011100_000000111111001000_000001111111100000_000000111111001000_000000000000011100_000000000000111100_000000000000111100_000000000000111100_000000000000111100_000000000000111100_000000000000111100_000000000000111100_000000000000011100_000000111111001000_000001111111100000_000000111111000000_000000000000000000_000000000000000000;
assign number[4] = 540'b000000000000000000_000000000000000000_000000000000000000_000100000000001000_001110000000011100_001111000000111100_001111000000111100_001111000000111100_001111000000111100_001111000000111100_001111000000111100_001111000000111100_001110000000011100_000100111111001000_000001111111100000_000000111111001000_000000000000011100_000000000000111100_000000000000111100_000000000000111100_000000000000111100_000000000000111100_000000000000111100_000000000000111100_000000000000011100_000000000000001000_000000000000000000_000000000000000000_000000000000000000_000000000000000000;
assign number[5] = 540'b000000000000000000_000000111111000000_000001111111100000_000100111111000000_001110000000000000_001111000000000000_001111000000000000_001111000000000000_001111000000000000_001111000000000000_001111000000000000_001111000000000000_001110000000000000_000100111111000000_000001111111100000_000000111111001000_000000000000011100_000000000000111100_000000000000111100_000000000000111100_000000000000111100_000000000000111100_000000000000111100_000000000000111100_000000000000011100_000000111111001000_000001111111100000_000000111111000000_000000000000000000_000000000000000000;
assign number[6] = 540'b000000000000000000_000000111111000000_000001111111100000_000100111111000000_001110000000000000_001111000000000000_001111000000000000_001111000000000000_001111000000000000_001111000000000000_001111000000000000_001111000000000000_001110000000000000_000100111111000000_000001111111100000_000100111111001000_001110000000011100_001111000000111100_001111000000111100_001111000000111100_001111000000111100_001111000000111100_001111000000111100_001111000000111100_001110000000011100_000100111111001000_000001111111100000_000000111111000000_000000000000000000_000000000000000000;
assign number[7] = 540'b000000000000000000_000000111111000000_000001111111100000_000000111111001000_000000000000011100_000000000000111100_000000000000111100_000000000000111100_000000000000111100_000000000000111100_000000000000111100_000000000000111100_000000000000011100_000000000000001000_000000000000000000_000000000000001000_000000000000011100_000000000000111100_000000000000111100_000000000000111100_000000000000111100_000000000000111100_000000000000111100_000000000000111100_000000000000011100_000000000000001000_000000000000000000_000000000000000000_000000000000000000_000000000000000000;
assign number[8] = 540'b000000000000000000_000000111111000000_000001111111100000_000100111111001000_001110000000011100_001111000000111100_001111000000111100_001111000000111100_001111000000111100_001111000000111100_001111000000111100_001111000000111100_001110000000011100_000100111111001000_000001111111100000_000100111111001000_001110000000011100_001111000000111100_001111000000111100_001111000000111100_001111000000111100_001111000000111100_001111000000111100_001111000000111100_001110000000011100_000100111111001000_000001111111100000_000000111111000000_000000000000000000_000000000000000000;
assign number[9] = 540'b000000000000000000_000000111111000000_000001111111100000_000100111111001000_001110000000011100_001111000000111100_001111000000111100_001111000000111100_001111000000111100_001111000000111100_001111000000111100_001111000000111100_001110000000011100_000100111111001000_000001111111100000_000000111111001000_000000000000011100_000000000000111100_000000000000111100_000000000000111100_000000000000111100_000000000000111100_000000000000111100_000000000000111100_000000000000011100_000000111111001000_000001111111100000_000000111111000000_000000000000000000_000000000000000000;


always @(*) begin

    index = (WIDTH*HEIGHT - ( (i_V_Cont-i_y)*WIDTH+(i_H_Cont-i_x)+1 ));

    // valid
    if (i_en && i_H_Cont-i_x >= 0 && i_H_Cont-i_x < WIDTH && i_V_Cont-i_y >= 0 && i_V_Cont-i_y < HEIGHT) begin
        case (i_speed)
            4'd0: begin o_valid = number[0][index]; end
            4'd1: begin o_valid = number[1][index]; end
            4'd2: begin o_valid = number[2][index]; end
            4'd3: begin o_valid = number[3][index]; end
            4'd4: begin o_valid = number[4][index]; end
            4'd5: begin o_valid = number[5][index]; end
            4'd6: begin o_valid = number[6][index]; end
            4'd7: begin o_valid = number[7][index]; end
            4'd8: begin o_valid = number[8][index]; end
            4'd9: begin o_valid = number[9][index]; end
            default: begin o_valid = 0; end
        endcase
    end else begin
        o_valid = 0;
    end
end

endmodule